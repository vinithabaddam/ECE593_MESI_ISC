/********************************************************************************
*
* Authors: Srijana Sapkota and Zeba Khan Rafi
* Reference: https://github.com/PrakashLuu/mesi_verification
* Reference: https://github.com/shruti2611/EE382M_project/blob/master/mesi_fifo/mesi_isc_define.v
* Reference: https://github.com/rdsalemi/uvmprimer/tree/master/16_Analysis_Ports_In_the_Testbench
* Reference: https://opencores.org/projects/mesi_isc
* Last Modified: March 6, 2019
*
* Description:	Driver for BFM. Inputs from tester are provided to
*				BFM's tasks through the FIFO.
********************************Change Log******************************************************* 
* Srijana S. and Zeba K. R.			3/6/2019			Created
********************************************************************************/

import mesi_isc_pkg::*;	
import uvm_pkg::*;
`include "uvm_macros.svh"

class driver extends uvm_component;
	`uvm_component_utils(driver)
	
	virtual mesi_isc_bfm bfm;
	
	uvm_get_port #(cpu_ip_s) cpu_ip_port;									  //declaring the get_port of the fifo
	
	
	function void build_phase(uvm_phase phase);
	
		if(!uvm_config_db #(virtual mesi_isc_bfm)::get(null, "*","bfm", bfm)) //extracting bfm handle from uvm db
			$fatal("Failed to get BFM");
		cpu_ip_port = new("cpu_ip_port",this);								  //instantiating the command fifo 
		
	endfunction : build_phase
	
	task run_phase(uvm_phase phase);
		  cpu_ip_s cpu_ip;													 //structure
		  
		  forever begin : command_loop
			 cpu_ip_port.get(cpu_ip);										 //pulling the cpu_ip structure(input to cpu) from fifo 
			 
			/* //check the cpu id to see which cpu to call 
			 if(cpu_ip.cpu_id == 'd3)
				bfm.send_ip_cpu3(cpu_ip);								     //calling bfm task to send commands to cpu 3
																			 //generated by the tester*/
			//just for now, change it to correct one
			bfm.send_ip_cpu(cpu_ip);

		  end : command_loop												  
	endtask : run_phase
	
	//constructor
	function new (string name, uvm_component parent);
		super.new(name, parent);
	endfunction : new
	
endclass: driver 
	
	
	
	
	
	
	
	
	